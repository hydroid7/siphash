module siphash;

endmodule